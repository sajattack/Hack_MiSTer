module Not16 (
    input [15:0] in,
    output wire [15:0] out
);

    _Not not0(in[0], out[0]);
    _Not not1(in[1], out[1]);
    _Not not2(in[2], out[2]);
    _Not not3(in[3], out[3]);
    _Not not4(in[4], out[4]);
    _Not not5(in[5], out[5]);
    _Not not6(in[6], out[6]);
    _Not not7(in[7], out[7]);
    _Not not8(in[8], out[8]);
    _Not not9(in[9], out[9]);
    _Not not10(in[10], out[10]);
    _Not not11(in[11], out[11]);
    _Not not12(in[12], out[12]);
    _Not not13(in[13], out[13]);
    _Not not14(in[14], out[14]);
    _Not not15(in[15], out[15]);


endmodule
