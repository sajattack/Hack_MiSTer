// nand2tetris Hack computer

module emu(
   //Master input clock
   input         CLK_50M,

   //Async reset from top-level module.
   //Can be used as initial reset.
   input         RESET,

   //Must be passed to hps_io module
   inout  [45:0] HPS_BUS,

   //Base video clock. Usually equals to CLK_SYS.
   output        CLK_VIDEO,

   //Multiple resolutions are supported using different CE_PIXEL rates.
   //Must be based on CLK_VIDEO
   output        CE_PIXEL,

   //Video aspect ratio for HDMI. Most retro systems have ratio 4:3.
   output  [7:0] VIDEO_ARX,
   output  [7:0] VIDEO_ARY,

   output  [7:0] VGA_R,
   output  [7:0] VGA_G,
   output  [7:0] VGA_B,
   output        VGA_HS,
   output        VGA_VS,
   output        VGA_DE,    // = ~(VBlank | HBlank)
   output        VGA_F1,
   output [1:0]  VGA_SL,

   output        LED_USER,  // 1 - ON, 0 - OFF.

   // b[1]: 0 - LED status is system status OR'd with b[0]
   //       1 - LED status is controled solely by b[0]
   // hint: supply 2'b00 to let the system control the LED.
   output  [1:0] LED_POWER,
   output  [1:0] LED_DISK,

   // I/O board button press simulation (active high)
   // b[1]: user button
   // b[0]: osd button
   output  [1:0] BUTTONS,

   output [15:0] AUDIO_L,
   output [15:0] AUDIO_R,
   output        AUDIO_S,   // 1 - signed audio samples, 0 - unsigned
   output  [1:0] AUDIO_MIX, // 0 - no mix, 1 - 25%, 2 - 50%, 3 - 100% (mono)

   //ADC
   inout   [3:0] ADC_BUS,

   //SD-SPI
   output        SD_SCK,
   output        SD_MOSI,
   input         SD_MISO,
   output        SD_CS,
   input         SD_CD,

   //High latency DDR3 RAM interface
   //Use for non-critical time purposes
   output        DDRAM_CLK,
   input         DDRAM_BUSY,
   output  [7:0] DDRAM_BURSTCNT,
   output [28:0] DDRAM_ADDR,
   input  [63:0] DDRAM_DOUT,
   input         DDRAM_DOUT_READY,
   output        DDRAM_RD,
   output [63:0] DDRAM_DIN,
   output  [7:0] DDRAM_BE,
   output        DDRAM_WE,

   //SDRAM interface with lower latency
   output        SDRAM_CLK,
   output        SDRAM_CKE,
   output [12:0] SDRAM_A,
   output  [1:0] SDRAM_BA,
   inout  [15:0] SDRAM_DQ,
   output        SDRAM_DQML,
   output        SDRAM_DQMH,
   output        SDRAM_nCS,
   output        SDRAM_nCAS,
   output        SDRAM_nRAS,
   output        SDRAM_nWE,

   input         UART_CTS,
   output        UART_RTS,
   input         UART_RXD,
   output        UART_TXD,
   output        UART_DTR,
   input         UART_DSR,

   // Open-drain User port.
   // 0 - D+/RX
   // 1 - D-/TX
   // 2..6 - USR2..USR6
   // Set USER_OUT to 1 to read from USER_IN.
   input   [6:0] USER_IN,
   output  [6:0] USER_OUT,

   input         OSD_STATUS
);


////////////////////////////  HPS I/O  //////////////////////////////////


`include "build_id.v"
parameter CONF_STR = {
   "Hack;;",
   "-;",
   "F,BIN;",
   "O1,Invert color,Yes,No;",
   "-;",
   "R0,Reset;",
   "V,v",`BUILD_DATE
};

wire  [1:0] buttons;
wire [31:0] status;

wire        ioctl_download;
wire [24:0] ioctl_addr;
wire [7:0] ioctl_dout;
wire        ioctl_wait;
wire        ioctl_wr;

hps_io #(.STRLEN($size(CONF_STR)>>3)) hps_io
(
   .clk_sys(clk_sys),
   .HPS_BUS(HPS_BUS),

   .conf_str(CONF_STR),

   .ioctl_download(ioctl_download),
   .ioctl_wr(ioctl_wr),
   .ioctl_addr(ioctl_addr),
   .ioctl_dout(ioctl_dout),
   .ioctl_wait(ioctl_wait),
   
   .buttons(buttons),
   .status(status),

   .ps2_key(ps2_key)
);


///////////////////////  CLOCK/RESET  ///////////////////////////////////

wire clock_locked;

wire clk_sys, clk_video;

pll pll
(
   .refclk(CLK_50M),
   .rst(0),
   .outclk_0(clk_sys),
   .outclk_1(clk_video),
   .locked(clock_locked)
);


wire reset = RESET | buttons[1] | status[0] | ioctl_download;

////////////////////////////  SYSTEM  ///////////////////////////////////
wire [14:0] addressM;
wire [15:0] outM, memOut, rom_out;
wire writeM;
wire [14:0] pc;
wire r, g, b, hsync, vsync;

CPU cpu(clk_sys, memOut, rom_out, reset, outM, writeM, addressM, pc);

assign CLK_VIDEO = clk_video;
assign VGA_R = {8{r^status[1]}};
assign VGA_G = {8{g^status[1]}};
assign VGA_B = {8{b^status[1]}};
assign VGA_HS = hsync;
assign VGA_VS = vsync;
assign VGA_DE = display_on;
assign VGA_SL = 0;
assign VGA_F1 = 0;
assign VIDEO_ARX = 8'd2;
assign VIDEO_ARY = 8'd1;
assign CE_PIXEL = 1'd1;

assign AUDIO_S = 0;

assign {UART_RTS, UART_TXD, UART_DTR} = 0;

assign {AUDIO_L, AUDIO_R} = 0;
assign AUDIO_S   = 0;
assign AUDIO_MIX = 0;

assign LED_USER  = 0;
assign LED_DISK  = ioctl_download;
assign LED_POWER = 0;
assign BUTTONS = 0;
assign ADC_BUS = 'Z;
assign USER_OUT = '1;
assign {SDRAM_DQ, SDRAM_A, SDRAM_BA, SDRAM_CKE, SDRAM_CLK, SDRAM_DQML, SDRAM_DQMH, SDRAM_nWE, SDRAM_nCAS, SDRAM_nRAS, SDRAM_nCS} = 'Z;
assign {DDRAM_CLK, DDRAM_BURSTCNT, DDRAM_ADDR, DDRAM_DIN, DDRAM_BE, DDRAM_RD, DDRAM_WE} = 0;
assign {SD_SCK, SD_MOSI, SD_CS} = 'Z;


////////////////////////////  INPUT  ////////////////////////////////////

wire [10:0] ps2_key;
wire [7:0] hack_scancode;

Keyboard keyboard(clk_sys, ps2_key, hack_scancode);

////////////////////////////  MEMORY & VIDEO ///////////////////////////////////  

reg count = 1'd0;
reg [15:0] rom_data_in = 16'd0;
reg [14:0] rom_addr_in = 15'd0;
reg rom_wr;

 dpram rom(
   .clock(clk_sys),
   .data(rom_data_in),
   .rdaddress(pc),
   .wraddress(rom_addr_in),
   .wren(rom_wr),
   .q(rom_out)
);
    
always @(posedge clk_sys) begin
   rom_wr <= 0;
   if (ioctl_wr) begin
      count <= count + 1'd1;
      if (count==0)
         rom_data_in[15:8] <= ioctl_dout;
      else begin
         rom_data_in[7:0] <= ioctl_dout;
         rom_addr_in <= ioctl_addr >> 1;
         rom_wr <= 1;
      end
   end else begin
      rom_addr_in <= rom_addr_in;
      count <= count;
      rom_data_in <= rom_data_in;
   end
end
 
 wire display_on;
 Memory mem(clk_sys, clk_video, reset, outM, writeM, addressM, memOut, hack_scancode, r, g, b, hsync, vsync, display_on);

endmodule
